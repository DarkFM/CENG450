----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:33:27 03/24/2017 
-- Design Name: 
-- Module Name:    sign_extend - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sign_extend is

    Port ( DISP_L : in  STD_LOGIC_VECTOR (8 downto 0);
           DISP_S : in  STD_LOGIC_VECTOR (5 downto 0);
           SEL : in  STD_LOGIC;
           EXTEND_OUT : out  STD_LOGIC_VECTOR (15 downto 0));
end sign_extend;

architecture Behavioral of sign_extend is

begin
--	process(DISP_L, DISP_S, SEL) begin
	
	EXTEND_OUT <=
			 std_logic_vector(resize(signed(DISP_L), EXTEND_OUT'length)) when SEL = '0' else
			 std_logic_vector(resize(signed(DISP_S), EXTEND_OUT'length));
--	end process;


end Behavioral;

